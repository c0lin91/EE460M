module DebounceAndSp(Button, DebouncedButton);

input Button;
output DebouncedButton;

endmodule
