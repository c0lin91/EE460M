//This module takes in the 4 digit BCD number and outputs the corresponding 7 segment LED values
module outputModule();

//stuff here

endmodule
