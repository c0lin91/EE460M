module inputModule(B0, B1, B2, B3, SW0, SW1, CLK, Q);

input B0, B1, B2, B3, SW0, SW1, CLK;
output [3:0] Q;

	

endmodule
